library verilog;
use verilog.vl_types.all;
entity colour_conversion is
end colour_conversion;
