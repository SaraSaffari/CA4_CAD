module colour_conversion();


endmodule 